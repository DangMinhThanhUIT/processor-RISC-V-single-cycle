`timescale 1ns/100ps
module Datapath_testbench();
reg CLK,  RegWrite, ALUSrc, MemWrite, MemRead, MemToReg;
reg [3:0] ALUControl;
reg [31:0] Instruction;
wire Sign, Zero;
initial begin
	#500 $stop;
end
initial begin
	RegWrite = 1'b1;
	ALUSrc = 0;
	ALUControl = 4'd0;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00010_00011_000_00001_0110011;
	#20// Add $1=$3+$2
	RegWrite = 1'b1;
	ALUSrc = 0;
	ALUControl = 4'd0;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00010_00011_000_00001_0110011;
	#20 // sub s4=s2-s3
	RegWrite = 1'b1;
	ALUSrc = 0;
	ALUControl = 4'd1;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b0100000_00011_00010_000_00100_0110011;
	#20 // or s5=s2|s3
	RegWrite = 1'b1;
	ALUSrc = 0;
	ALUControl = 4'd3;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00011_00010_110_00101_0110011;
	#20 // and s6=s2&s3
	RegWrite = 1'b1;
	ALUSrc = 0;
	ALUControl = 4'd2;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00011_00010_111_00110_0110011;
	#20 // sll s7=s2<<s3
	RegWrite = 1'b1;
	ALUSrc = 0;
	ALUControl = 4'd4;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00011_00010_001_00111_0110011;
	#20 // slt s8 = (s2 << s3) ? 1:0
	RegWrite = 1'b1;
	ALUSrc = 0;
	ALUControl = 4'd5;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00011_00010_010_01000_0110011;
	#20 // addi s9 = s2 + 20
	RegWrite = 1'b1;
	ALUSrc = 1;
	ALUControl = 4'd0;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b000000010100_00010_000_01001_0010011;
	#20 // xori s10=s2^20
	RegWrite = 1'b1;
	ALUSrc = 1;
	ALUControl = 4'd6;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b000000010100_00010_100_01010_0010011;
	#20 // ori s11=s2|20
 	RegWrite = 1'b1;
	ALUSrc = 1;
	ALUControl = 4'd3;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b000000010100_00010_110_01011_0010011;
	#20 // andi s12=s2&20
	RegWrite = 1'b1;
	ALUSrc = 1;
	ALUControl = 4'd2;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b000000010100_00010_111_01100_0010011;
	#40 // sw M[s2+20]=s1
   RegWrite = 1'b0;
	ALUSrc = 1;
	ALUControl = 4'd0;
	MemWrite = 1'b1;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00001_00010_010_10100_0100011;
	#40 // lw s14=M[s2+20]
	RegWrite = 1'b1;
	ALUSrc = 1;
	ALUControl = 4'd0;
	MemWrite = 1'b0;
	MemRead = 1'b1;
	MemToReg = 1'b1;
	Instruction = 32'b000000010100_00010_010_01110_0000011 ;
	#40 // xor s15=s2^s3
	RegWrite = 1'b1;
	ALUSrc = 0;
	ALUControl = 4'd6;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00011_00010_100_01111_0110011;
	#40 // srl s16=s2>>s3
	RegWrite = 1'b1;
	ALUSrc = 0;
	ALUControl = 4'd7;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00011_00010_101_10000_0110011;
	#20 // sltu s17=s2<s3 ? 1:0
	RegWrite = 1'b1;
	ALUSrc = 0;
	ALUControl = 4'd8;
	MemWrite = 1'b0;
	MemRead = 1'b0;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00011_00010_011_10001_0110011;
	#20 // slli s18=s2<< 2
	RegWrite = 1'b1;
	ALUSrc = 1;
	ALUControl = 4'd4;
	MemWrite = 1'b0;
	MemRead = 1'b1;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00010_00010_001_10010_0010011 ;
	#20// srli s19=s2>> 2
	RegWrite = 1'b1;
	ALUSrc = 1;
	ALUControl = 4'd7;
	MemWrite = 1'b0;
	MemRead = 1'b1;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_00010_00010_001_10011_0010011 ;
	#20// slti s20=s2<20 ? 1:0
	RegWrite = 1'b1;
	ALUSrc = 1;
	ALUControl = 4'd5;
	MemWrite = 1'b0;
	MemRead = 1'b1;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_10100_00010_010_10100_0010011 ;
	#20// sltiu s21=s2< 20 ?1:0
	RegWrite = 1'b1;
	ALUSrc = 1;
	ALUControl = 4'd8;
	MemWrite = 1'b0;
	MemRead = 1'b1;
	MemToReg = 1'b0;
	Instruction = 32'b0000000_10100_00010_010_10101_0010011 ;
	#20// lui $22=20<<12
	RegWrite = 1'b1;
	ALUSrc = 1;
	ALUControl = 4'd4;
	MemWrite = 1'b0;
	MemRead = 1'b1;
	MemToReg = 1'b0;
	Instruction = 32'b00000000000000010100_10110_0110111 ;
end
Datapath Datapath1(.CLK(CLK),.RegWrite (RegWrite),.ALUSrc (ALUSrc),.ALUControl (ALUControl),. MemWrite(MemWrite),. MemRead(MemRead),
. MemToReg(MemToReg),.Instruction (Instruction),. Sign(Sign),.Zero (Zero));
initial
begin
	CLK = 0;
	forever #10 CLK=~CLK;
end
endmodule