module Adder(input [31:0] a, b, output [31:0] y);
	assign y = $signed(a) + $signed(b);
endmodule